module deboucner(
);
