`timescale 1ns / 1ps

module ssd_driver(
    input clk,
    input [3:0] disp1,    // in order from left to right
    input [3:0] disp2,
    input [3:0] disp3,
    input [3:0] disp4,
    input [0:0] blink,
    output reg [7:0] cathodes,
    output reg [3:0] anodes
);

endmodule
